--
-- Definition of a single port ROM for KCPSM3 program defined by uclock.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity uclock is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end uclock;
--
architecture low_level_definition of uclock is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "0D0000A4E00CE00BE00AE009E008E007E006E005E004E003E002E001E0000000";
attribute INIT_01 of ram_1024_x_18  : label is "40490091501200ED50374041501E40545012400D0091012000C30115C0010C00";
attribute INIT_02 of ram_1024_x_18  : label is "5812006D541C4020401200A8542C400D0091541C40450091541C404D0091541C";
attribute INIT_03 of ram_1024_x_18  : label is "541C40520091541C40410091541C404C0091401200A8E005E004E408E507E606";
attribute INIT_04 of ram_1024_x_18  : label is "5812006DC1015055404F0091541C4020401200AC5448400D0091541C404D0091";
attribute INIT_05 of ram_1024_x_18  : label is "401200ACE00CC002600C541C400D00915460404E0091401200ACE40BE50AE609";
attribute INIT_06 of ram_1024_x_18  : label is "1620588B01EC401200AC00A4E00C0000541C400D0091541C40460091541C4046";
attribute INIT_07 of ram_1024_x_18  : label is "009181011420588B01EC548B403A009181011520588B01EC548B403A00918101";
attribute INIT_08 of ram_1024_x_18  : label is "000E0001013400E70125A000000E00005C8B443C5C8B453C5C8B4618548B400D";
attribute INIT_09 of ram_1024_x_18  : label is "50A220024000A000009D4F0140950185549A20104000A000810101E27010A000";
attribute INIT_0A of ram_1024_x_18  : label is "013D00BC01600E09A00000BC01600E06A000C000A001600CA000CF01409D0185";
attribute INIT_0B of ram_1024_x_18  : label is "4F0D009D7F100120A0000148A000014E50BA2002A000015350B62001600C00E7";
attribute INIT_0C of ram_1024_x_18  : label is "810150D34F08B0004F0DFF10009554DB2008400082101210012040BD8101B000";
attribute INIT_0D of ram_1024_x_18  : label is "400000E400FAEF2000E440C3012240C600EA00E758D94120C10100EA54C65120";
attribute INIT_0E of ram_1024_x_18  : label is "0F79009D0F53A000009D0F08A000009D0F20A000009D0F0D40DF4F01B0002010";
attribute INIT_0F of ram_1024_x_18  : label is "009D0F65009D0F76009D0F4F410A009D0F78009D0F61009D0F74009D0F6E009D";
attribute INIT_10 of ram_1024_x_18  : label is "009D009D0F72009D0F4500E7009D0F77009D0F6F009D0F6C009D0F66009D0F72";
attribute INIT_11 of ram_1024_x_18  : label is "009D0F4D009D0F53009D0F50009D0F43009D0F4B00E4A000009D0F72009D0F6F";
attribute INIT_12 of ram_1024_x_18  : label is "0F69009D0F6C009D0F61009D0F76009D0F6E009D0F49A000009D0F3E009D0F33";
attribute INIT_13 of ram_1024_x_18  : label is "0F6C009D0F41A000009D0F65009D0F6D009D0F69009D0F54A000009D0F64009D";
attribute INIT_14 of ram_1024_x_18  : label is "009D0F4FA000009D009D0F46009D0F4FA000009D0F6D009D0F72009D0F61009D";
attribute INIT_15 of ram_1024_x_18  : label is "A000009D0F65009D0F76009D0F69009D0F74009D0F63009D0F41A000009D0F4E";
attribute INIT_16 of ram_1024_x_18  : label is "F0208201F120017E70E08E018201F020003A8201F0208201F120017E70E00220";
attribute INIT_17 of ram_1024_x_18  : label is "81010130A000F020000D8201F0208201F120017E70E08E018201F020003A8201";
attribute INIT_18 of ram_1024_x_18  : label is "EC01ED00C00063016200E515E414E313E212E111E010A000803AC1015D7FC00A";
attribute INIT_19 of ram_1024_x_18  : label is "82E8419A8001599FE303C2E80000B350924063036202F530D42065016400C001";
attribute INIT_1A of ram_1024_x_18  : label is "E204A30382E841AF800159ADE303C2E80000A300920063056204E303E202A303";
attribute INIT_1B of ram_1024_x_18  : label is "010041C9E10751BF413C81016107E108010041C9E10851B7413C91006108E305";
attribute INIT_1C of ram_1024_x_18  : label is "5010610A600755DB501061096006E106010041C9E10651C7411881016106E107";
attribute INIT_1D of ram_1024_x_18  : label is "6414631362126111601000A4E00CC00151DB2002600C55DB5010610B600855DB";
attribute INIT_1E of ram_1024_x_18  : label is "1200B80001E87010A000C0F6B80080C6A000A0DFBC00407BB8004061A0006515";
attribute INIT_1F of ram_1024_x_18  : label is "000000000000000000000000A0009200B80001E8701081010206920002060206";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "43FC8001AC008D01000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "D3F74FDD3FF8DF7DF837DFEAF77DFDF7DF7DFEAAFDFDF7DF7FDDDCFC3AAAAAA8";
attribute INITP_01 of ram_1024_x_18 : label is "CCCF333332CB2CC93EFFFD7D766F443670BBDBD3FCBCA0AFD2CFD2728FE8DDDD";
attribute INITP_02 of ram_1024_x_18 : label is "4A19B1619B1619B0B333332CCBCCB33332CCCCB3333332CCCCCCCECCF33CCCCC";
attribute INITP_03 of ram_1024_x_18 : label is "0009B19A2C9989980038D34343423B523B523B529775142977514143AC2AAA5D";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "F500000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"0D0000A4E00CE00BE00AE009E008E007E006E005E004E003E002E001E0000000",
                INIT_01 => X"40490091501200ED50374041501E40545012400D0091012000C30115C0010C00",
                INIT_02 => X"5812006D541C4020401200A8542C400D0091541C40450091541C404D0091541C",
                INIT_03 => X"541C40520091541C40410091541C404C0091401200A8E005E004E408E507E606",
                INIT_04 => X"5812006DC1015055404F0091541C4020401200AC5448400D0091541C404D0091",
                INIT_05 => X"401200ACE00CC002600C541C400D00915460404E0091401200ACE40BE50AE609",
                INIT_06 => X"1620588B01EC401200AC00A4E00C0000541C400D0091541C40460091541C4046",
                INIT_07 => X"009181011420588B01EC548B403A009181011520588B01EC548B403A00918101",
                INIT_08 => X"000E0001013400E70125A000000E00005C8B443C5C8B453C5C8B4618548B400D",
                INIT_09 => X"50A220024000A000009D4F0140950185549A20104000A000810101E27010A000",
                INIT_0A => X"013D00BC01600E09A00000BC01600E06A000C000A001600CA000CF01409D0185",
                INIT_0B => X"4F0D009D7F100120A0000148A000014E50BA2002A000015350B62001600C00E7",
                INIT_0C => X"810150D34F08B0004F0DFF10009554DB2008400082101210012040BD8101B000",
                INIT_0D => X"400000E400FAEF2000E440C3012240C600EA00E758D94120C10100EA54C65120",
                INIT_0E => X"0F79009D0F53A000009D0F08A000009D0F20A000009D0F0D40DF4F01B0002010",
                INIT_0F => X"009D0F65009D0F76009D0F4F410A009D0F78009D0F61009D0F74009D0F6E009D",
                INIT_10 => X"009D009D0F72009D0F4500E7009D0F77009D0F6F009D0F6C009D0F66009D0F72",
                INIT_11 => X"009D0F4D009D0F53009D0F50009D0F43009D0F4B00E4A000009D0F72009D0F6F",
                INIT_12 => X"0F69009D0F6C009D0F61009D0F76009D0F6E009D0F49A000009D0F3E009D0F33",
                INIT_13 => X"0F6C009D0F41A000009D0F65009D0F6D009D0F69009D0F54A000009D0F64009D",
                INIT_14 => X"009D0F4FA000009D009D0F46009D0F4FA000009D0F6D009D0F72009D0F61009D",
                INIT_15 => X"A000009D0F65009D0F76009D0F69009D0F74009D0F63009D0F41A000009D0F4E",
                INIT_16 => X"F0208201F120017E70E08E018201F020003A8201F0208201F120017E70E00220",
                INIT_17 => X"81010130A000F020000D8201F0208201F120017E70E08E018201F020003A8201",
                INIT_18 => X"EC01ED00C00063016200E515E414E313E212E111E010A000803AC1015D7FC00A",
                INIT_19 => X"82E8419A8001599FE303C2E80000B350924063036202F530D42065016400C001",
                INIT_1A => X"E204A30382E841AF800159ADE303C2E80000A300920063056204E303E202A303",
                INIT_1B => X"010041C9E10751BF413C81016107E108010041C9E10851B7413C91006108E305",
                INIT_1C => X"5010610A600755DB501061096006E106010041C9E10651C7411881016106E107",
                INIT_1D => X"6414631362126111601000A4E00CC00151DB2002600C55DB5010610B600855DB",
                INIT_1E => X"1200B80001E87010A000C0F6B80080C6A000A0DFBC00407BB8004061A0006515",
                INIT_1F => X"000000000000000000000000A0009200B80001E8701081010206920002060206",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"43FC8001AC008D01000000000000000000000000000000000000000000000000",    
               INITP_00 => X"D3F74FDD3FF8DF7DF837DFEAF77DFDF7DF7DFEAAFDFDF7DF7FDDDCFC3AAAAAA8",
               INITP_01 => X"CCCF333332CB2CC93EFFFD7D766F443670BBDBD3FCBCA0AFD2CFD2728FE8DDDD",
               INITP_02 => X"4A19B1619B1619B0B333332CCBCCB33332CCCCB3333332CCCCCCCECCF33CCCCC",
               INITP_03 => X"0009B19A2C9989980038D34343423B523B523B529775142977514143AC2AAA5D",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"F500000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE uclock.vhd
--
------------------------------------------------------------------------------------
